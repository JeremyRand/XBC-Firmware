# ====================================================================
#
#      hal_m68k_mcf52xx_mcf5272_mcf5272c3.cdl
#
#      Motorola mcf5272c3 evaluation board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================

cdl_package CYGPKG_HAL_M68K_MCF52xx_MCF5272_MCF5272C3 {
    display         "Motorola mcf5272c3 evaluation board"
    parent          CYGPKG_HAL_M68K_MCF52xx_MCF5272
    define_header   hal_m68k_mcf52xx_mcf5272_mcf5272c3.h
    include_dir     cyg/hal

    description   "The  Motorola  mcf5272c3  evaluation  board  platform   HAL
                package should be used when targeting the actual hardware  for
                the Motorola mcf5272c3 evaluation board platform."

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_m68k_mcf52xx_mcf5272.h>"
    }

    compile     plf_startup.c hal_diag.c

#    implements      CYGINT_HAL_DEBUG_GDB_STUBS
#    implements      CYGINT_HAL_DEBUG_GDB_STUBS_BREAK

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_m68k.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H <pkgconf/hal_m68k_mcf52xx_mcf5272.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_m68k_mcf52xx_mcf5272_mcf5272c3.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display         "Startup type"
        flavor          data
        legal_values    {"RAM" "ROM"}
        default_value   {"RAM"}
	    no_define
	    define -file system.h CYG_HAL_STARTUP

        description   "When targeting the Motorola mcf5272c3 evaluation  board
                    it is expected that the image will be downloaded into  RAM
                    via the Motorola dBUG monitor."

    }

    cdl_option CYGHWR_HAL_SYSTEM_CLOCK_MHZ {
       display          "System clock speed in MHz"
       flavor data
       legal_values     66
       default_value    66

       description    "This  option  identifies  the  system  clock  that  the
                    processor uses.  This value is used to set clock  dividers
                    for some devices."

    }

    cdl_option CYGHWR_HAL_M68K_MCF52xx_MCF5272_MCF5272C3_DIAG_BAUD {
       display          "Diagnostic Serial Port Baud Rate"
       flavor data
       legal_values     9600 19200 38400 115200
       default_value    9600

       description    "This  option  selects  the  baud  rate  used  for   the
                    diagnostic port.  Note: this should match the value chosen
                    for the GDB port if  the diagnostic and  GDB port are  the
                    same."

    }

    cdl_option CYGHWR_HAL_M68K_MCF52xx_MCF5272_MCF5272C3_GDB_BAUD {
       display          "GDB Serial Port Baud Rate"
       flavor data
       legal_values     9600 19200 38400 115200
       default_value    9600

       description    "This option controls  the baud  rate used  for the  GDB
                    connection."

    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none

        description   "Set the periodic timer  on  the  mcf5272  to  1  ms  or
                    1000000 ns."

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    1000
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    1000000
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE

        description   "Global build  options including  control over  compiler
                    flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "m68k-elf" }

            description       "This option specifies  the command prefix  used
                            when invoking the build tools."

        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-m5200 -malign-int -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-thunks=3 -finit-priority -fomit-frame-pointer" }
            description       "This option controls the global compiler  flags
                            which are used to compile all packages by default.
                            Individual  packages  may  define  options   which
                            override these global flags."

        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-m5200 -g -nostdlib -Wl,--gc-sections -Wl,-static" }

            description       "This option controls  the global linker  flags.
                            Individual  packages  may  define  options   which
                            override these global flags."

        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define

            description       "This option enables the  building  of  the  GDB
                            stubs for the  board.   The  common  HAL  controls
                            takes care of most of  the build process, but  the
                            final conversion from ELF image to binary data  is
                            handled by the  platform CDL, allowing  relocation
                            of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.srec : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O srec $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "m68k_mcf52xx_mcf5272_mcf5272c3_ram" : \
	                                        "m68k_mcf52xx_mcf5272_mcf5272c3_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_m68k_mcf52xx_mcf5272_mcf5272c3_ram.ldi>" : \
                                                    "<pkgconf/mlt_m68k_mcf52xx_mcf5272_mcf5272c3_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_m68k_mcf52xx_mcf5272_mcf5272c3_ram.h>" : \
                                                    "<pkgconf/mlt_m68k_mcf52xx_mcf5272_mcf5272c3_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        requires      { CYG_HAL_STARTUP == "RAM" }
        parent        CYGPKG_HAL_ROM_MONITOR

        description       "Support  can  be  enabled  for  boot  ROMs  or  ROM
                        monitors  which  contain  GDB  stubs.   This   support
                        changes various eCos semantics such as the encoding of
                        diagnostic output,  and  the  overriding  of  hardware
                        interrupt vectors."

    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }

        description       "Enable this option if this program is to be used as
                        a ROM monitor, i.e.  applications will be loaded  into
                        RAM on the  board, and  this ROM  monitor may  process
                        exceptions   or   interrupts   generated   from    the
                        application.  This enables features such as  utilizing
                        a  separate  interrupt   stack  when  exceptions   are
                        generated."

    }
}
