# ====================================================================
#
#      wallclock.cdl
#
#      eCos wallclock configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  nickg
# Contributors:
# Date:           1999-07-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_WALLCLOCK {
    display       "Wallclock device"
    include_dir   cyg/io

    define_header wallclock.h
    description   "
        The wallclock device provides real time stamps, as opposed
        to the eCos kernel timers which typically just count the
        number of clock ticks since the hardware was powered up.
        Depending on the target platform this device may involve
        interacting with a suitable clock chip, or it may be
        emulated by using the kernel timers."

    compile       wallclock.cxx

    cdl_interface CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS {
        display       "Number of wallclock hardware implementations"
        no_define
    }

    cdl_interface CYGINT_WALLCLOCK_IMPLEMENTATIONS {
        display       "Number of wallclock implementations"
        no_define
        requires      1 == CYGINT_WALLCLOCK_IMPLEMENTATIONS
    }

    cdl_interface CYGINT_WALLCLOCK_SET_GET_MODE_SUPPORTED {
        display       "Wallclock driver supports set/get mode"
        no_define
    }

    cdl_option CYGSEM_WALLCLOCK_MODE {
        display       "Wallclock mode"
        flavor        data
        legal_values  { "init_get" "set_get" }
        default_value { CYGINT_WALLCLOCK_SET_GET_MODE_SUPPORTED ? \
                        "set_get" : "init_get" }
        requires      { CYGINT_WALLCLOCK_SET_GET_MODE_SUPPORTED || \
                        CYGSEM_WALLCLOCK_MODE == "init_get" }
        no_define
        description   "
            The wallclock driver can be used in one of two
            modes. Set/get mode allows time to be kept during power
            off (assuming there's a battery backed clock). Init/get
            mode is slightly smaller and can be used when there is no
            battery backed clock - in this mode time 0 is the time of
            the board power up."
    }

    cdl_option CYGSEM_WALLCLOCK_SET_GET_MODE {
        display     "Wallclock set/get mode"
        calculated  { CYGSEM_WALLCLOCK_MODE == "set_get" ? 1 : 0 }
    }

    cdl_component CYGPKG_IO_WALLCLOCK_IMPLEMENTATION {
        display "Wallclock implementation"
        flavor none
        no_define
        description "Implementations of the wallclock device."

        cdl_option CYGPKG_WALLCLOCK_EMULATE {
            default_value { 0 == CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS }
            display       "Wallclock emulator"
            implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
            compile       emulate.cxx
            requires      CYGPKG_KERNEL
            define_proc {
                puts $::cdl_header "#undef CYGSEM_WALLCLOCK_SET_GET_MODE"
            }
            description   "
                When this option is enabled, a wallclock device will be
                emulated using the kernel real-time clock."
        }

        cdl_option CYGIMP_WALLCLOCK_NONE {
            display       "No wallclock"
            default_value { !CYGPKG_KERNEL && 0 == CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS }
            implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
            description   "Disables the wallclock."
        }
    }

    cdl_component CYGPKG_IO_WALLCLOCK_OPTIONS {
        display "Wallclock build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_WALLCLOCK_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_WALLCLOCK_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_IO_WALLCLOCK_TESTS {
            display "Wallclock tests"
            flavor  data
            no_define
            calculated { CYGPKG_KERNEL ? "tests/wallclock tests/wallclock2" : "" }
            description   "
                This option specifies the set of tests for the
                wallclock device."
        }
    }
}
