# ====================================================================
#
#      mfc_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for MCF5272
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================

cdl_package CYGPKG_NET_MCF5272_ETH_DRIVERS {
    display       "MCF5272 ethernet driver"
    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0
    implements    CYGHWR_NET_DRIVERS
    include_dir   cyg/devs/eth
    description   "MCF5272 Ethernet driver"
    compile       -library=libextras.a if_mcf5272.c nbuf.c

    cdl_component CYGPKG_NET_MCF5272_ETH_DRIVERS_OPTIONS {
        display "MCF5272 ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_NET_MCF5272_ETH_DRIVERS_RX_NUM_BDS {
                display       "The number of receive buffer descriptors"
                flavor        data
                legal_values  2 to 2048
                default_value 256
                description   "
                    This option specifies the number of buffer descriptors that
                    the driver should allocated for the receive side."
            }

        cdl_option CYGPKG_NET_MCF5272_ETH_DRIVERS_TX_NUM_BDS {
                display       "The number of transmit buffer descriptors"
                flavor        data
                legal_values  2 to 2048
                default_value 128
                description   "
                    This option specifies the number of buffer descriptors that
                    the driver should allocated for the transmit side."
            }


        cdl_option CYGPKG_NET_MCF5272_ETH_DRIVERS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the MCF5272 ethernet driver package. These flags are used in addition
                to the set of global flags."
        }
    }
}
