# ====================================================================
#
#      mn10300_asb2305_eth.cdl
#
#      Ethernet drivers - support for AMD PCnet ethernet controller
#      on the ASB2305 board.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      dhowells
# Contributors:   jskov
# Date:           2001-07-23
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_MN10300_ASB2305 {
    display       "MN10300 ASB2305 board ethernet driver"
    description   "Ethernet driver for MN10300 ASB2305 onboard ethernet device."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_MN10300_AM33_ASB2305

    include_dir   cyg/io

    # FIXME: This really belongs in the AMD_PCNET package
    cdl_interface CYGINT_DEVS_ETH_AMD_PCNET_REQUIRED {
        display   "AMD PCNET ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_AMD_PCNET_INL <cyg/io/mn10300_asb2305_eth.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_AMD_PCNET_CFG <pkgconf/devs_eth_mn10300_asb2305.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component CYGPKG_DEVS_ETH_MN10300_ASB2305_ETH0 {
        display       "ASB2305 ethernet port 0 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the ethernet device driver for the
            ASB2305 port 0."

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_AMD_PCNET_REQUIRED

        cdl_option CYGNUM_DEVS_ETH_MN10300_ASB2305_ETH0_RX_RING_SIZE {
            display       "Size of RX ring for ETH0"
            flavor        data
            default_value 4
            legal_values  { 4 8 16 32 64 128 }
            description   "
                This option sets the size of the RX ring."
        }

        cdl_option CYGNUM_DEVS_ETH_MN10300_ASB2305_ETH0_TX_RING_SIZE {
            display       "Size of TX ring for ETH0"
            flavor        data
            default_value 16
            legal_values  { 4 8 16 32 64 128 }
            description   "
                This option sets the size of the TX ring."
        }

        cdl_option CYGDAT_DEVS_ETH_MN10300_ASB2305_ETH0_NAME {
            display       "Device name for the ETH0 ethernet port 0 driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device for the
                ASB2305 port 0."
        }

        cdl_component CYGSEM_DEVS_ETH_MN10300_ASB2305_ETH0_SET_ESA {
            display       "Set the ethernet station address"
            flavor        bool
            default_value 0
            description   "Enabling this option will allow the ethernet
            station address to be forced to the value set by the
            configuration.  This may be required if the hardware does
            not include a serial EEPROM for the ESA."
            
            cdl_option CYGDAT_DEVS_ETH_MN10300_ASB2305_ETH0_ESA {
                display       "The ethernet station address"
                flavor        data
                default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
                description   "The ethernet station address"
            }
        }
    }
}
