# ====================================================================
#
#      flash_iq80310.cdl
#
#      FLASH memory - Hardware support on Cyclone IQ80310
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  msalter
# Contributors:
# Date:           2000-10-10
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_IQ80310 {
    display       "Cyclone IQ80310 FLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  CYGPKG_HAL_ARM_IQ80310

    implements    CYGHWR_IO_FLASH_DEVICE
    implements    CYGHWR_IO_FLASH_DEVICE_NOT_IN_RAM
    implements    CYGHWR_IO_FLASH_BLOCK_LOCKING

    include_dir   .
    include_files ; # none _exported_ whatsoever
    description   "FLASH memory device support for Cyclone IQ80310"
    compile       iq80310_flash.c

    make -priority 1 {
        flash_erase_block.o: $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        echo " .globl flash_erase_block_end" >>flash_erase_block.s
        echo "flash_erase_block_end:" >>flash_erase_block.s
        $(CC) $(CFLAGS) -c -o flash_erase_block.o flash_erase_block.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_erase_block.o
    }
    make -priority 1 {
        flash_program_buf.o: $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        echo " .globl flash_program_buf_end" >>flash_program_buf.s
        echo "flash_program_buf_end:" >>flash_program_buf.s
        $(CC) $(CFLAGS) -c -o flash_program_buf.o flash_program_buf.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_program_buf.o
    }
    make -priority 1 {
        flash_query.o: $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        echo " .globl flash_query_end" >>flash_query.s
        echo "flash_query_end:" >>flash_query.s
        $(CC) $(CFLAGS) -c -o flash_query.o flash_query.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_query.o
    }
    make -priority 1 {
        flash_lock_block.o: $(REPOSITORY)/$(PACKAGE)/src/flash_lock_block.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_lock_block.c
        echo " .globl flash_lock_block_end" >>flash_lock_block.s
        echo "flash_lock_block_end:" >>flash_lock_block.s
        $(CC) $(CFLAGS) -c -o flash_lock_block.o flash_lock_block.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_lock_block.o
    }
    make -priority 1 {
        flash_unlock_block.o: $(REPOSITORY)/$(PACKAGE)/src/flash_unlock_block.c
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_unlock_block.c
        echo " .globl flash_unlock_block_end" >>flash_unlock_block.s
        echo "flash_unlock_block_end:" >>flash_unlock_block.s
        $(CC) $(CFLAGS) -c -o flash_unlock_block.o flash_unlock_block.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_unlock_block.o
    }
}

