# ====================================================================
#
#      frv400_eth_drivers.cdl
#
#      Ethernet drivers - support for i82559 ethernet controller
#      on the Fujitsu FR-V400
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov, hmt, gthomas
# Date:           2001-02-28
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_FRV_FRV400 {
    display       "FRV400 ethernet driver"
    description   "
	Ethernet drivers for Fujitsu FR-V400 board."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_PCI
    requires      CYGPKG_DEVS_ETH_NS_DP83902A

    implements    CYGHWR_NET_DRIVER_ETH0
    include_dir   cyg/io

#    compile       -library=libextras.a if_frv400.c

    # FIXME: This really belongs in the NS DP83902A package
    cdl_interface CYGINT_DEVS_ETH_NS_DP83902A_REQUIRED {
        display   "NS DP83902A ethernet driver required"
    }
	
    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NS_DP83902A_INL <cyg/io/devs_eth_frv400.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NS_DP83902A_CFG <pkgconf/devs_eth_frv_frv400.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component CYGPKG_DEVS_ETH_FRV400_ETH0 {
        display       "CF ethernet port driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the ethernet device driver for a
            CF card."

        implements CYGINT_DEVS_ETH_NS_DP83902A_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_FRV400_ETH0_NAME {
            display       "Device name for the ETH0 ethernet driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device."
        }

        cdl_component CYGSEM_DEVS_ETH_FRV400_ETH0_SET_ESA {
            display       "Set the ethernet station address"
            flavor        bool
            default_value 0
            description   "Enabling this option will allow the ethernet
            station address to be forced to the value set by the
            configuration.  This may be required if the hardware does
            not include a serial EEPROM for the ESA."
            
            cdl_option CYGDAT_DEVS_ETH_FRV400_ETH0_ESA {
                display       "The ethernet station address"
                flavor        data
                default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
                description   "The ethernet station address"
            }
        }
    }

    cdl_component CYGPKG_DEVS_ETH_FRV400_OPTIONS {
        display "PCMCIA ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_FRV400_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the PCMCIA ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }
}

# EOF frv400_eth_drivers.cdl
