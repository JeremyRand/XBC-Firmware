# ====================================================================
#
#      hal_arm_aeb.cdl
#
#      AEB1 board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  gthomas
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_AEB {
    display       "ARM AEB-1 evaluation board"
    parent        CYGPKG_HAL_ARM
    requires      ! CYGHWR_THUMB
    define_header hal_arm_aeb.h
    include_dir   cyg/hal
    hardware
    description   "
        The aeb HAL package provides the support needed to run
        eCos on a ARM AEB-1 eval board."

    compile       hal_diag.c aeb_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_ARM_ARCH_ARM7
    implements    CYGINT_HAL_TESTS_NO_CACHES

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_aeb.h>"

        puts $::cdl_header "#define CYGPRI_KERNEL_TESTS_DHRYSTONE_PASSES 100000"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the AEB-1 eval board it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using onboard
            debug software such as Angel or eCos GDB stubs.  Select 'rom'
            when building a stand-alone application which will be put
            into ROM."
    }


    cdl_option CYGHWR_HAL_ARM_AEB_REVISION {
        display       "AEB board revision"
        flavor        data
        default_value {"B"}
        legal_values  {"B" "C"}
        description   "
            The AEB-1 eval board exists in two revisions. Revision B
            has 128kB of memory and a flawed CPU which means caches
            must be disabled. Revision C has 256kB of memory and can
            run with caches enabled."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The AEB board has only one serial port. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The AEB board has only one serial port.  This option
            chooses which port will be used for diagnostic output."
     }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    (240000/16)
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm7di -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm7di -Wl,--gc-sections -Wl,-static -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires ! CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. This is a bit convoluted as it involves prepending
                the image with a special header used by the AEB firmware
                to keep track of multiple ROM images. This header includes
                a checksum making it necessary to build twice."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PACKAGE>/src/gdb_module.c
                @sh -c "mkdir -p src $(dir $@)"
                # First build version with no checksum.
                $(CC) -c $(INCLUDE_PATH) -Wp,-MD,deps.tmp -I$(dir $<) $(CFLAGS) -o src/gdb_module_ncs.o $<
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o src/gdb_module_ncs.tmp src/gdb_module_ncs.o
                $(OBJCOPY) --strip-debug --change-addresses=0xFBFF4000 src/gdb_module_ncs.tmp src/gdb_module_ncs.img
                $(OBJCOPY) -O binary src/gdb_module_ncs.img src/gdb_module_ncs.bin
                @rm src/gdb_module_ncs.tmp src/gdb_module_ncs.img
                # Prepare dependency file
                @echo $@ ": \\" > $(notdir $@).deps
                @echo $(wildcard $(PREFIX)/lib/*) " \\" >> $(notdir $@).deps
                @tail +2 deps.tmp >> $(notdir $@).deps
                @echo >> $(notdir $@).deps
                @rm deps.tmp
                # Then build version with checksum from previously built image.
                @cp $(dir $<)flash_cksum.tcl src/
                $(CC) -c -DCHECKSUM=`src/flash_cksum.tcl src/gdb_module_ncs.bin` $(INCLUDE_PATH) -I$(dir $<) $(CFLAGS) -o src/gdb_module.o $<
                $(CC) $(LDFLAGS) -L$(PREFIX)/lib -Ttarget.ld -o src/gdb_module.tmp src/gdb_module.o
                $(OBJCOPY) --strip-debug --change-addresses=0xFBFF4000 src/gdb_module.tmp $(@:.bin=.img)
                $(OBJCOPY) -O binary $(@:.bin=.img) src/gdb_module.bin
                uuencode src/gdb_module.bin gdb_module.bin | tr '`' ' ' > $(@:.bin=.img.UU)
                @rm src/gdb_module.tmp src/gdb_module_ncs.bin
		@mv src/gdb_module.bin $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { (CYGHWR_HAL_ARM_AEB_REVISION == "B" &&           \
                      CYG_HAL_STARTUP == "RAM") ? "arm_aeb_ram" :     \
                     (CYGHWR_HAL_ARM_AEB_REVISION == "B" &&           \
                      CYG_HAL_STARTUP == "ROM") ? "arm_aeb_rom" :     \
                     (CYGHWR_HAL_ARM_AEB_REVISION == "C" &&           \
                      CYG_HAL_STARTUP == "RAM") ? "arm_aebC_ram" :    \
                      "arm_aebC_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { (CYGHWR_HAL_ARM_AEB_REVISION == "B" &&           \
                          CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_aeb_ram.ldi>" :     \
                         (CYGHWR_HAL_ARM_AEB_REVISION == "B" &&           \
                          CYG_HAL_STARTUP == "ROM") ? "<pkgconf/mlt_arm_aeb_rom.ldi>" :     \
                         (CYGHWR_HAL_ARM_AEB_REVISION == "C" &&           \
                          CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_aebC_ram.ldi>" :    \
                         "<pkgconf/mlt_arm_aebC_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { (CYGHWR_HAL_ARM_AEB_REVISION == "B" &&           \
                          CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_aeb_ram.h>" :     \
                         (CYGHWR_HAL_ARM_AEB_REVISION == "B" &&           \
                          CYG_HAL_STARTUP == "ROM") ? "<pkgconf/mlt_arm_aeb_rom.h>" :     \
                         (CYGHWR_HAL_ARM_AEB_REVISION == "C" &&           \
                          CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_arm_aebC_ram.h>" :    \
                          "<pkgconf/mlt_arm_aebC_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }
}
