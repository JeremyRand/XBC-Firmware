# ====================================================================
#
#      hal_calm16_ceb.cdl
#
#      CalmRISC16 Core Eval Board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  bartv
# Contributors:
# Date:           2001-02-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_CALM16_CEB {
    display  "CalmRISC16 core evaluation board"
    parent        CYGPKG_HAL_CALM16
    include_dir   cyg/hal
    description   "
           The Core eval board HAL package should be used when targetting the
           actual hardware."

    compile       hal_diag.c platform.S plf_misc.c ser.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT_GUARANTEED

    cdl_option CYGBLD_HAL_TARGET_H {
        display       "Variant header"
        flavor        data
	no_define
	calculated { "<pkgconf/hal_calm16_core.h>" }
	define -file system.h CYGBLD_HAL_TARGET_H
        description   "Variant header."

        define_proc {
            puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_calm16_ceb.h>"
            puts $::cdl_system_header ""
            puts $::cdl_system_header "/* Make sure we get the CORE type definitions for HAL_PLATFORM_CPU */"
            puts $::cdl_system_header "#include CYGBLD_HAL_TARGET_H"
	    puts $::cdl_system_header "#define HAL_PLATFORM_BOARD    \"Ceb\""
	    puts $::cdl_system_header "#define HAL_PLATFORM_EXTRA    \"\""
	    puts $::cdl_system_header ""
        }
				      
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM"}
        default_value {"ROM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
            Currently only ROM startup type is supported."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  57600
        default_value 57600
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  57600
        default_value 57600
        description   "
            This option controls the baud rate used for the GDB connection."
    }

    cdl_option CYGBLD_BUILD_GDB_STUBS {
	display "Build GDB stub ROM image"
	default_value 0
	parent CYGBLD_GLOBAL_OPTIONS
	requires { CYG_HAL_STARTUP == "ROM" }
	requires CYGSEM_HAL_ROM_MONITOR
	requires CYGBLD_BUILD_COMMON_GDB_STUBS
	requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
	requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
	requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
	requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
	requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
	no_define
	description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

	make -priority 320 {
	    <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
	    $(OBJCOPY) -O binary $< $@
	}
    }


    cdl_option CYGNUM_HAL_BREAKPOINT_LIST_SIZE {
        display       "Number of breakpoints supported by the HAL."
        flavor        data
        default_value 25
        description   "
            This option determines the number of breakpoints supported by the HAL."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The Atlas board has only one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The Atlas board has only one serial port.  This option
           chooses which port will be used for diagnostic output."
     }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "calm16_ceb_ram" : \
                                                "calm16_ceb_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_calm16_ceb_ram.ldi>" : \
                                                    "<pkgconf/mlt_calm16_ceb_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_calm16_ceb_ram.h>" : \
                                                    "<pkgconf/mlt_calm16_ceb_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "Generic" "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "Generic" : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        description   "
            Support can be enabled for three different varieties of ROM monitor.
            This support changes various eCos semantics such as the encoding
            of diagnostic output, or the overriding of hardware interrupt
            vectors.
            Firstly there is \"Generic\" support which prevents the HAL
            from overriding the hardware vectors that it does not use, to
            instead allow an installed ROM monitor to handle them. This is
            the most basic support which is likely to be common to most
            implementations of ROM monitor.
            \"CygMon\" provides support for the Cygnus ROM Monitor.
            And finally, \"GDB_stubs\" provides support when GDB stubs are
            included in the ROM monitor or boot ROM."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 1
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."
    
        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            compile -library=libextras.a
    
            make -priority 325 {
                <PREFIX>/bin/redboot.srec : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-all $< $(@:.srec=.img)
                $(OBJCOPY) -O srec $< $@
            }
        }
    }

}
